`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:44:06 12/30/2019 
// Design Name: 
// Module Name:    reg_bank 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module reg_bank(
input [3:0] op1,
input [3:0] op2,
output reg[15:0] op1_out,
output reg[15:0] op2_out,
input clk
    );

reg [3:0] temp1;
reg [3:0] temp2;
always @(posedge clk)
begin
case (temp1)
4'b0000: op1_out [15:0] =16'b0000000000001000;
4'b0001: op1_out [15:0] =16'b0000000000001000;
4'b0010: op1_out [15:0] =16'b0000000000001000;
4'b0011: op1_out [15:0] =16'b0000000000001000;
4'b0100: op1_out [15:0] =16'b0000000000000000;
4'b0101: op1_out [15:0] =16'b0000000000000000;
4'b0110: op1_out [15:0] =16'b0000000000000000;
4'b0111: op1_out [15:0] =16'b0000000000000000;
4'b1000: op1_out [15:0] =16'b0000000000000000;
4'b1001: op1_out [15:0] =16'b0000000000000000;
4'b1010: op1_out [15:0] =16'b0000000000000000;
4'b1011: op1_out [15:0] =16'b0000000000000000;
4'b1100: op1_out [15:0] =16'b0000000000000000;
4'b1101: op1_out [15:0] =16'b0000000000000000;
4'b1110: op1_out [15:0] =16'b0000000000000000;
4'b1111: op1_out [15:0] =16'b0000000000000000;
endcase

case (temp2)
4'b0000: op2_out [15:0] =16'b0000000000111000;
4'b0001: op2_out [15:0] =16'b0000000000111000;
4'b0010: op2_out [15:0] =16'b0000000000000000;
4'b0011: op2_out [15:0] =16'b0000000000000000;
4'b0100: op2_out [15:0] =16'b0000000000000000;
4'b0101: op2_out [15:0] =16'b0000000000000000;
4'b0110: op2_out [15:0] =16'b0000000000000000;
4'b0111: op2_out [15:0] =16'b0000000000000000;
4'b1000: op2_out [15:0] =16'b0000000000000000;
4'b1001: op2_out [15:0] =16'b0000000000000000;
4'b1010: op2_out [15:0] =16'b0000000000000000;
4'b1011: op2_out [15:0] =16'b0000000000000000;
4'b1100: op2_out [15:0] =16'b0000000000000000;
4'b1101: op2_out [15:0] =16'b0000000000000000;
4'b1110: op2_out [15:0] =16'b0000000000000000;
4'b1111: op2_out [15:0] =16'b0000000000000000;
endcase
end
endmodule
